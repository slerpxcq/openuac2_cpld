`timescale 1ns/1ps

module tb_dop_detector;
endmodule